library IEEE;

use IEEE.std_logic_1164.all;
use work.user_defines.all;

entity generate_fsm_tb is
end entity;
