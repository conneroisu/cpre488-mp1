-- library declaration
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
-- entity
entity ppm_generation is
	port (
	);
end ppm_generation;

architecture arc of ppm_generation is
begin
end arc;
