library IEEE;

-- Blank for now

use IEEE.std_logic_1164.all;
use work.user_defines.all;

entity detect_fsm_tb is
end entity;